* IRLZ44N switching Peltier with 12V supply (low-side switching)

* PWM gate signal (500 kHz, 50% duty)
VG GPIO 0 PULSE(0 3.3 0 130n 130n 1u 2u); *130ns is the max propogation delay from the SN74HC245 datasheet

* Gate
RG GPIO G_p 33
RPULL G_p 0 100k
Vprobe G G_p 0

* 12V Power Supply
VDD vdd 0 DC 12

* Peltier Load
VPelt vdd Peltier 0
RPelt Peltier D 2
CPelt D 0 1p

* MOSFET
X1 D G 0 irlz44n

* Simulation control
.tran 0.1u 2u

.control
run
plot V(D) V(G) 
plot I(VPelt) 
plot I(Vprobe)
.endc



* Inline IRLZ44N model
.SUBCKT irlz44n 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=2.08819 LAMBDA=0.0038193 KP=67.9211
+CGSO=1.59143e-05 CGDO=3.04562e-08
RS 8 3 0.014066
D1 3 1 MD
.MODEL MD D IS=4.4574e-09 RS=0.007275 N=1.40246 BV=55
+IBV=0.00025 EG=1.14011 XTI=3.00078 TT=0
+CJO=8.92434e-10 VJ=4.94724 M=0.75496 FC=0.5
RDS 3 1 2.2e+06
RD 9 1 0.00179971
RG 2 7 2.4114
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.15401e-09 VJ=0.859156 M=0.642548 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.64838e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS